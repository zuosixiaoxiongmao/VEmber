module core

pub struct Vec {
	x f32
	y f32
}

pub struct Vec3 {
	x f32
	y f32
	z f32
}

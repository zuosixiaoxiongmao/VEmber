module core

pub struct Object {

}
module gate

import core {Entity, System, ServicerComponent}
import parts {ConfigComponent}

pub struct GateComponet {

}
module utilities

